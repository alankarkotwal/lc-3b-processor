//`include "misc/mux.v"
//`include "misc/demux.v"

module controller();

endmodule