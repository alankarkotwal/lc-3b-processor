// Skeleton file for the LC-3b processor

`include "alu/alu.v"
`include "reg-file/register_file.v"

module lc_3b();

endmodule
