// Skeleton file for the LC-3b processor

`include "datapath.v"
`include "controller.v"

module lc_3b();

endmodule
