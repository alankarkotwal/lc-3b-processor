`include "reg-file/register_file.v"
`include "alu/alu.v"

module datapath();

endmodule